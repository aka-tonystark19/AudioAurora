
module fft_acc (
	clk_clk,
	lights_readdata,
	reset_reset_n);	

	input		clk_clk;
	output	[8:0]	lights_readdata;
	input		reset_reset_n;
endmodule
