
module fft_acc (
	clk_clk,
	reset_reset_n,
	lights_readdata);	

	input		clk_clk;
	input		reset_reset_n;
	output	[8:0]	lights_readdata;
endmodule
